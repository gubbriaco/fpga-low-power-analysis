library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library work;
use work.MyDefinitions.all;


entity TopArchitectureTB is
end TopArchitectureTB;




architecture Behavioral of TopArchitectureTB is

	-- System Signal definitions
	signal i_clk : std_logic := '0';
	constant T_CLK : Time := 10 ns;
	signal i_rst : std_logic := '0';

	-- Components declaration
	component TopArchitecture is
		port (
			a, b, c, d : in std_logic_vector(nBitsInputs-1 downto 0);
			sel1, sel2 : in std_logic_vector(nBitsSels-1 downto 0);
			clk, rst : in std_logic;
			z : out std_logic_vector(nBitsInputs downto 0)
		);
	end component;
	
	-- TopArchitecture Signals definitions
	signal aTB : std_logic_vector(nBitsInputs-1 downto 0) := (others=>'0');
	signal bTB : std_logic_vector(nBitsInputs-1 downto 0) := (others=>'0');
	signal cTB : std_logic_vector(nBitsInputs-1 downto 0) := (others=>'0');
	signal dTB : std_logic_vector(nBitsInputs-1 downto 0) := (others=>'0');
	signal sel1TB : std_logic_vector(nBitsSels-1 downto 0) := (others=>'0');
	signal sel2TB : std_logic_vector(nBitsSels-1 downto 0) := (others=>'0');
	signal zTB : std_logic_vector(nBitsInputs downto 0);
	

	begin
	
		uut : TopArchitecture port map(
				aTB,
				bTB,
				cTB,
				dTB,
				sel1TB,
				sel2TB,
				i_clk,
				i_rst,
				zTB
			);
		
		
		clk_process : process
        begin
				wait for T_CLK/2;
          i_clk <= not i_clk;
     end process clk_process;
	 
		-- rst_process : process
        -- begin
				-- wait for 20ns;
           -- i_rst <= not i_rst;
				-- wait for 10ns;
				-- i_rst <= not i_rst;
     -- end process rst_process;
	 
	 
		uut_process : process
			begin
				wait for 100ns;
				i_rst <= '1';
				wait for 10ns;
				i_rst <= '0';
			
aTB <= "01001011000010011011010100001101";
bTB <= "11111110001011101001001100111111";
cTB <= "00110110111001101111101010101111";
dTB <= "00110111010000100011101011011101";
sel1TB <= "01011011";
sel2TB <= "11001100";
wait for T_CLK;
aTB <= "11100001000110110011001011000011";
bTB <= "01010010110001011000100101100110";
cTB <= "11100000100011010010010010110010";
dTB <= "00101100100010011011000100110001";
sel1TB <= "10110001";
sel2TB <= "11101010";
wait for T_CLK;
aTB <= "00001100111111100011100101010011";
bTB <= "11111101001001000111001011001010";
cTB <= "00011100001110001101000011000100";
dTB <= "10101010010110000101000111011111";
sel1TB <= "11011101";
sel2TB <= "00010100";
wait for T_CLK;
aTB <= "00011001101001011101110010101100";
bTB <= "10000111100101011000111011111000";
cTB <= "01011101110010000101001100010000";
dTB <= "10000100111101010011001110000111";
sel1TB <= "01010111";
sel2TB <= "01111000";
wait for T_CLK;
aTB <= "00011101011100111111101010001100";
bTB <= "11001110001110110100011101011111";
cTB <= "00101100110011000100001001110001";
dTB <= "01111101001101111001100011111001";
sel1TB <= "10100000";
sel2TB <= "10101111";
wait for T_CLK;
aTB <= "10000001010011100100100100000101";
bTB <= "00010101000001001011111001100110";
cTB <= "00000110001111000111000001011101";
dTB <= "01110111110100110010110110111100";
sel1TB <= "01001101";
sel2TB <= "11000000";
wait for T_CLK;
aTB <= "10100001011010011010000010000001";
bTB <= "00111010000111001011100111111011";
cTB <= "00011001101111111001011101101000";
dTB <= "01011011000110111000001101111100";
sel1TB <= "00101011";
sel2TB <= "11110010";
wait for T_CLK;
aTB <= "01111100100111101001011001111010";
bTB <= "11100111011001010110010100001100";
cTB <= "01111001101010011110110011000111";
dTB <= "10001011110111000110110101010101";
sel1TB <= "00110111";
sel2TB <= "10010011";
wait for T_CLK;
aTB <= "01101110101110101001001100000110";
bTB <= "11001101000000111101010011001100";
cTB <= "00110011101000000101010010100101";
dTB <= "10101010011001111001010011101111";
sel1TB <= "00100111";
sel2TB <= "01100110";
wait for T_CLK;
aTB <= "00101000001101011101000101101001";
bTB <= "01111000111101111101011101010011";
cTB <= "01001111011000001110001100010000";
dTB <= "11111110100110110101100010111100";
sel1TB <= "01110011";
sel2TB <= "10001101";
wait for T_CLK;
aTB <= "01001000000100110010111111000110";
bTB <= "11110000110111111010010001101110";
cTB <= "01000110111100110000010001111111";
dTB <= "11001011001101101010100010101101";
sel1TB <= "00110011";
sel2TB <= "01000100";
wait for T_CLK;
aTB <= "10110110010000100100011000010010";
bTB <= "11110111111111111101011000000111";
cTB <= "00111001010000010001000100000000";
dTB <= "11100100110101010011000111000100";
sel1TB <= "11100110";
sel2TB <= "10100000";
wait for T_CLK;
aTB <= "10101011000100110000100000001000";
bTB <= "00111000001001000111011010101101";
cTB <= "00110000100000110111100100001100";
dTB <= "01000011000001110100100110001100";
sel1TB <= "01001001";
sel2TB <= "11011100";
wait for T_CLK;
aTB <= "01011000110110010010110011011110";
bTB <= "00110111100110101100001001100111";
cTB <= "11011011001101001010010010001101";
dTB <= "01110011001101010000010101000110";
sel1TB <= "10001101";
sel2TB <= "10010101";
wait for T_CLK;
aTB <= "00100010011001011011000101110011";
bTB <= "00101010010110100100010000011000";
cTB <= "00101101011110111001111010000101";
dTB <= "01111111001001000101001011010000";
sel1TB <= "10011001";
sel2TB <= "01000000";
wait for T_CLK;
aTB <= "10000001011111000010001110110110";
bTB <= "10111010101011000100110101101010";
cTB <= "00100011011101100010000001111001";
dTB <= "10010100001011001001001110011001";
sel1TB <= "00111101";
sel2TB <= "11011001";
wait for T_CLK;
aTB <= "00111010000111000111101101110011";
bTB <= "01001001110110011110001101100110";
cTB <= "00001001101110010101011001111100";
dTB <= "00100011000010001010100011110010";
sel1TB <= "01000010";
sel2TB <= "11110000";
wait for T_CLK;
aTB <= "11000100011110000010010011001100";
bTB <= "11001101101011101011000101010000";
cTB <= "11100011000010111110011100111001";
dTB <= "00100011011011001000100110001110";
sel1TB <= "01100010";
sel2TB <= "10011110";
wait for T_CLK;
aTB <= "01001001101011111100110101110100";
bTB <= "01000001100111110000101001111100";
cTB <= "11101100100100011101010001111011";
dTB <= "01001000001110100100010000011000";
sel1TB <= "00000111";
sel2TB <= "11000011";
wait for T_CLK;
aTB <= "01000000101001101110011110100110";
bTB <= "11011100111010100110011001110101";
cTB <= "00111100011110001000100001101101";
dTB <= "11100010101010000000110000000000";
sel1TB <= "10001101";
sel2TB <= "00001011";
wait for T_CLK;
aTB <= "00010011001001011011010000000010";
bTB <= "01100100101000011010011101111111";
cTB <= "01100011000101000001100110011110";
dTB <= "01111011001101101111111010011000";
sel1TB <= "01110111";
sel2TB <= "11101101";
wait for T_CLK;
aTB <= "00011010100111101011011110011101";
bTB <= "11000000001111111111100111011001";
cTB <= "11110011001101110001101111111111";
dTB <= "11001111011110111000111010100001";
sel1TB <= "10110101";
sel2TB <= "11101000";
wait for T_CLK;
aTB <= "01100000111000000100010000110110";
bTB <= "10100110000100011100001100000010";
cTB <= "11111100000100100111111100011000";
dTB <= "10101110011110010111010110100110";
sel1TB <= "11010110";
sel2TB <= "10011110";
wait for T_CLK;
aTB <= "11000101010001011010110101111011";
bTB <= "10100100111110000011010011101101";
cTB <= "00010001100100100011111101100100";
dTB <= "01100001010101101001010111101000";
sel1TB <= "10000100";
sel2TB <= "01011110";
wait for T_CLK;
aTB <= "00000011000001011101011100101111";
bTB <= "00100101111000011101001000010101";
cTB <= "00000100100110001010010011010111";
dTB <= "11001010000111100000110010010101";
sel1TB <= "00000011";
sel2TB <= "10111000";
wait for T_CLK;
aTB <= "10110111011001010000100100001000";
bTB <= "10011110110101101110001100011011";
cTB <= "11101101101010000001000010110100";
dTB <= "11000000001000111100001001100010";
sel1TB <= "10001001";
sel2TB <= "01101101";
wait for T_CLK;
aTB <= "11111100000100011110110111001000";
bTB <= "01110011001101001111110101011000";
cTB <= "10110111001111011101101100011011";
dTB <= "10101011000000000000010001111001";
sel1TB <= "10101000";
sel2TB <= "00110000";
wait for T_CLK;
aTB <= "01011010000000011111110110100010";
bTB <= "00100110101000001111000000111000";
cTB <= "11111110101001100101111100011111";
dTB <= "00110101001001000111101011011101";
sel1TB <= "11010101";
sel2TB <= "00011101";
wait for T_CLK;
aTB <= "10101001100001000100110111011011";
bTB <= "11000111111110111111101100101011";
cTB <= "11001110111001010010101101110101";
dTB <= "11000101101000011111101010000011";
sel1TB <= "11110001";
sel2TB <= "11111011";
wait for T_CLK;
aTB <= "00000100110100011011000110110000";
bTB <= "10110001101100100000010101100110";
cTB <= "11011010111001100111100010111110";
dTB <= "11010110100000011010111100101011";
sel1TB <= "00001100";
sel2TB <= "00000101";
wait for T_CLK;
aTB <= "10000110111001001110100101101011";
bTB <= "11101100000000000011010101010101";
cTB <= "11100011111111100000111110011101";
dTB <= "01001110111100111001011001100011";
sel1TB <= "01100100";
sel2TB <= "11100100";
wait for T_CLK;
aTB <= "11111101011011100101111110011001";
bTB <= "11111001001011001000001111011000";
cTB <= "11010010110101100110010111010101";
dTB <= "01011101110100101010011010100011";
sel1TB <= "01010111";
sel2TB <= "01100100";
wait for T_CLK;
aTB <= "10100110001101010011100110101011";
bTB <= "00001100001110011011100001100000";
cTB <= "11111001011100010000001111101100";
dTB <= "00110000010011110101000110010100";
sel1TB <= "00000110";
sel2TB <= "00011111";
wait for T_CLK;
aTB <= "00000110101110101111111111010100";
bTB <= "11000111000001011000010011101110";
cTB <= "10111111100101000010111011011110";
dTB <= "10100011010001111101010011000000";
sel1TB <= "11010110";
sel2TB <= "00001110";
wait for T_CLK;
aTB <= "10111000101101010110111001100110";
bTB <= "11110100101110111111110010010101";
cTB <= "10000111111110100110111010000110";
dTB <= "10110010010001001111000000100100";
sel1TB <= "01011010";
sel2TB <= "00110101";
wait for T_CLK;
aTB <= "10100110101110010101001110011110";
bTB <= "10100111111011000100100011101000";
cTB <= "11100100100011011110001010001100";
dTB <= "00010111010110000100110101111010";
sel1TB <= "00110001";
sel2TB <= "10011101";
wait for T_CLK;
aTB <= "00100111111101110110011000011010";
bTB <= "00001011011101010111010111011111";
cTB <= "10101110000110110000001010011011";
dTB <= "00111010000000101101101100110110";
sel1TB <= "00110101";
sel2TB <= "00110010";
wait for T_CLK;
aTB <= "10111010101010100000110011000100";
bTB <= "11000001111000101011000001110111";
cTB <= "11001100000101101101100111000001";
dTB <= "01100101110110100110100111110010";
sel1TB <= "01010001";
sel2TB <= "00011111";
wait for T_CLK;
aTB <= "11000011010011110011111010111000";
bTB <= "10000100100101100101010100001011";
cTB <= "01111111110110010001111010010111";
dTB <= "10101111100010000111111000101110";
sel1TB <= "10010001";
sel2TB <= "11011011";
wait for T_CLK;
aTB <= "11011100101011001100010100000000";
bTB <= "00000010000001100011011011011001";
cTB <= "10011011001100100010000011111010";
dTB <= "00100110011010111000110001111111";
sel1TB <= "00011011";
sel2TB <= "00001100";
wait for T_CLK;
aTB <= "11111010101001111111111010001000";
bTB <= "11110111111000011010100111101110";
cTB <= "10011011010010001100000000000010";
dTB <= "01110010010111001001110000100001";
sel1TB <= "01111010";
sel2TB <= "01000000";
wait for T_CLK;
aTB <= "00000100101010100110101101001100";
bTB <= "11001110000110010001110111110101";
cTB <= "10101001010000110010000010000101";
dTB <= "10100011111010000010111111010001";
sel1TB <= "10110001";
sel2TB <= "11100110";
wait for T_CLK;
aTB <= "11110000100011111000110101111100";
bTB <= "10111110000001101010101100100101";
cTB <= "00010000101011011100010111111010";
dTB <= "00111110011011110100001010011001";
sel1TB <= "01010101";
sel2TB <= "10101001";
wait for T_CLK;
aTB <= "10001111000010011101101100001110";
bTB <= "01101010001010010110010000101000";
cTB <= "00101100010100010111001010110001";
dTB <= "01110011000000101100001110011001";
sel1TB <= "01000101";
sel2TB <= "00111010";
wait for T_CLK;
aTB <= "01111011001011010011100110100100";
bTB <= "00110111101010000100100001001100";
cTB <= "10011111000000001100010111000011";
dTB <= "00100010010111000101110011111111";
sel1TB <= "00110111";
sel2TB <= "11111001";
wait for T_CLK;
aTB <= "11111111010010101010101101101010";
bTB <= "01100110101110001011101111100011";
cTB <= "01010101000010001101011100100000";
dTB <= "11000010001000010000100001010010";
sel1TB <= "01101011";
sel2TB <= "10100011";
wait for T_CLK;
aTB <= "01010000100000000110111101011101";
bTB <= "01110101101100001011100010000101";
cTB <= "11100001111110011010011010111001";
dTB <= "01000110011001011100010111011111";
sel1TB <= "00101100";
sel2TB <= "00000001";
wait for T_CLK;
aTB <= "11111110100010101100011001110010";
bTB <= "01000111000110001110001001101001";
cTB <= "11011101100110010110100101100010";
dTB <= "01010011000101100111011101101010";
sel1TB <= "11010011";
sel2TB <= "10011001";
wait for T_CLK;
aTB <= "10001011010101111100110000000001";
bTB <= "00001110000011110101011100000001";
cTB <= "11101110011111010011101010000111";
dTB <= "01010100010000111011101011010011";
sel1TB <= "11010111";
sel2TB <= "10100000";
wait for T_CLK;
aTB <= "01111000111010100100101010101110";
bTB <= "10110100101100100100001111011100";
cTB <= "10001101000001111001111111101101";
dTB <= "11011011110101111110001010111000";
sel1TB <= "10001000";
sel2TB <= "01101001";
wait for T_CLK;
aTB <= "01100111101010101110110000000001";
bTB <= "10001110110101110010011100101100";
cTB <= "00110010100001010101101111100001";
dTB <= "10011010010010001101101010000000";
sel1TB <= "10011101";
sel2TB <= "01010001";
wait for T_CLK;
aTB <= "11000111101010000000010110001011";
bTB <= "00110001011010000001011110011000";
cTB <= "00110100110001001101010000101001";
dTB <= "10110001110111011010101111111000";
sel1TB <= "01011011";
sel2TB <= "00000000";
wait for T_CLK;
aTB <= "01101001101111100001001110011010";
bTB <= "11101000011011000011010111111011";
cTB <= "00000111011111010010111011000111";
dTB <= "11011000101110001000010110100010";
sel1TB <= "11100110";
sel2TB <= "00101100";
wait for T_CLK;
aTB <= "10010100100100001110011011110010";
bTB <= "10001000000001000000010001110001";
cTB <= "10001111100011000011001111001011";
dTB <= "10001111010100101000000100100101";
sel1TB <= "00100001";
sel2TB <= "00001001";
wait for T_CLK;
aTB <= "11111101101101100011000101111111";
bTB <= "00000011000010101010111001010100";
cTB <= "10111101100100111011001000110010";
dTB <= "11011100111111101010000101101111";
sel1TB <= "11101001";
sel2TB <= "01010010";
wait for T_CLK;
aTB <= "00010000000000001100010101001100";
bTB <= "10011000010010010110101110100001";
cTB <= "01101011000010001011000011000011";
dTB <= "10001010101010010001001010100100";
sel1TB <= "00001001";
sel2TB <= "11101000";
wait for T_CLK;
aTB <= "01001010100011011001110011011100";
bTB <= "11011111101100100001010010010100";
cTB <= "00100110000010011111000101000100";
dTB <= "00011101010101011100101011100100";
sel1TB <= "00101100";
sel2TB <= "10001011";
wait for T_CLK;
aTB <= "11101100000111000000001111101001";
bTB <= "11111100001110111111001110000000";
cTB <= "10110001110010011111101110100000";
dTB <= "11001001100100111111011011101011";
sel1TB <= "00001101";
sel2TB <= "00110101";
wait for T_CLK;
aTB <= "01101011011010110111011000011110";
bTB <= "10111100101101011011001111001101";
cTB <= "01011001011111110001001001100100";
dTB <= "11011100001000010110001101001111";
sel1TB <= "11110001";
sel2TB <= "11010000";
wait for T_CLK;
aTB <= "00111010100010010001011000101101";
bTB <= "10010110110101111001000110110000";
cTB <= "10010101100110000000000001100100";
dTB <= "00110100101011101111111000011010";
sel1TB <= "11110101";
sel2TB <= "10111100";
wait for T_CLK;
aTB <= "11111011111110000100000100100111";
bTB <= "01110000011100101000100100110011";
cTB <= "11011001011000001010110000110101";
dTB <= "10001000000110101101101010001110";
sel1TB <= "11111111";
sel2TB <= "00011011";
wait for T_CLK;
aTB <= "10100110100111000101011011110100";
bTB <= "11111111011111001011101111010110";
cTB <= "11101011111101111100111000100010";
dTB <= "10101001101011010111110000001100";
sel1TB <= "01001000";
sel2TB <= "10000000";
wait for T_CLK;
aTB <= "01110010000011111101001011001000";
bTB <= "10001001100001101101011111101100";
cTB <= "11011000111010010001001110100000";
dTB <= "10101000111101001110110000111110";
sel1TB <= "10101011";
sel2TB <= "11110100";
wait for T_CLK;
aTB <= "01110111000010110011000101001011";
bTB <= "10001000100101010010000110011100";
cTB <= "01000011101001010011010100111001";
dTB <= "10101001011100010110110001100011";
sel1TB <= "01011100";
sel2TB <= "00101100";
wait for T_CLK;
aTB <= "11011100110101010010010110110101";
bTB <= "11001011000110011000111011110001";
cTB <= "10101000101100101111001010100001";
dTB <= "11111011011011000011010110000100";
sel1TB <= "11010010";
sel2TB <= "11110010";
wait for T_CLK;
aTB <= "01101110001010000100010110000011";
bTB <= "01110110000000010011101110101101";
cTB <= "01111111111100110110011111111010";
dTB <= "10111000101001100010001000000011";
sel1TB <= "01101011";
sel2TB <= "10100011";
wait for T_CLK;
aTB <= "10001011100100111101001001111111";
bTB <= "11000111100000110110101100010000";
cTB <= "10100011001101100010100100101000";
dTB <= "10000110100010010000010010111000";
sel1TB <= "01111100";
sel2TB <= "00000001";
wait for T_CLK;
aTB <= "00011110110111011100000010000101";
bTB <= "01001100001111101010000110011100";
cTB <= "00001001110100001010111000011000";
dTB <= "00000100000010010001100011110011";
sel1TB <= "01010010";
sel2TB <= "11101001";
wait for T_CLK;
aTB <= "01011111010000100010101010111000";
bTB <= "00000111100000111001001110110111";
cTB <= "11100110100011000000101111100111";
dTB <= "01010011000010011110001111011010";
sel1TB <= "00000000";
sel2TB <= "00100000";
wait for T_CLK;
aTB <= "11011000101101011000111110100001";
bTB <= "00001010111010000000101101011000";
cTB <= "10111100101001001100000011000011";
dTB <= "10011100001111111100011100000111";
sel1TB <= "01001010";
sel2TB <= "00110011";
wait for T_CLK;
aTB <= "00100010001111010001100011001010";
bTB <= "01100010110111001011000111011110";
cTB <= "10001100000010110101011101101011";
dTB <= "00110110111000000000001011011100";
sel1TB <= "01010110";
sel2TB <= "10110011";
wait for T_CLK;
aTB <= "10011000000011111100101100000011";
bTB <= "00011010010000101100111000111110";
cTB <= "00100100110011101110100001001000";
dTB <= "00100000101010000110001101000110";
sel1TB <= "00000110";
sel2TB <= "00101101";
wait for T_CLK;
aTB <= "10011110001110000111010111101111";
bTB <= "11101100110101110010111111101001";
cTB <= "11111111000010101001000100101101";
dTB <= "01010001000010011011000100000100";
sel1TB <= "00111111";
sel2TB <= "10000101";
wait for T_CLK;
aTB <= "01001111001010010101101011010001";
bTB <= "00000101010100011101000101100110";
cTB <= "10101101000111110000000100001111";
dTB <= "11110001010011000001111010111011";
sel1TB <= "01100100";
sel2TB <= "10101010";
wait for T_CLK;
aTB <= "00100001001010000000011011111110";
bTB <= "11110111000001100000011101100101";
cTB <= "01001100110100011011110110011001";
dTB <= "01101111100111101000100010010010";
sel1TB <= "11001011";
sel2TB <= "01000101";
wait for T_CLK;
aTB <= "10000111010000001001010001000100";
bTB <= "00111001011010011100001001001010";
cTB <= "11100100010110000111101100110101";
dTB <= "10011110110010001110100100101101";
sel1TB <= "00100101";
sel2TB <= "10111000";
wait for T_CLK;
aTB <= "11011000001000110010000011010000";
bTB <= "00110101100110010111100000001011";
cTB <= "10110100110111001001100111010111";
dTB <= "00101110010101110001110010000011";
sel1TB <= "10000111";
sel2TB <= "01111111";
wait for T_CLK;
aTB <= "00110011100100100111011010010010";
bTB <= "11111000011001011010110111010000";
cTB <= "01101001100010110101100011110111";
dTB <= "00100101100000100101100011001010";
sel1TB <= "01010001";
sel2TB <= "01011001";
wait for T_CLK;
aTB <= "10111001000110110001101111110000";
bTB <= "01010111000001111110011001011100";
cTB <= "00001101101010100000001100000101";
dTB <= "11101000011110001010000101111000";
sel1TB <= "01100111";
sel2TB <= "01001001";
wait for T_CLK;
aTB <= "00111101101001000000011101011101";
bTB <= "01000111001000100011110110100100";
cTB <= "00111110010111101110011010100101";
dTB <= "00001000100110000111000110111010";
sel1TB <= "10110000";
sel2TB <= "10001100";
wait for T_CLK;
aTB <= "10100000001111000000100011010101";
bTB <= "00000011001110000111101011110101";
cTB <= "10100010100110000000111001110001";
dTB <= "10000000011010000010100010001000";
sel1TB <= "00010001";
sel2TB <= "01100101";
wait for T_CLK;
aTB <= "01110011001110010000100101001110";
bTB <= "10101111101111101101111111110100";
cTB <= "00110010111111111000001111111011";
dTB <= "11001010000101011011001110000111";
sel1TB <= "11100011";
sel2TB <= "10000001";
wait for T_CLK;
aTB <= "00110110110010111010110101000110";
bTB <= "01010101100001111111011100010000";
cTB <= "01101000100101110101001100110011";
dTB <= "01011101101010101000010111101001";
sel1TB <= "10011011";
sel2TB <= "00011101";
wait for T_CLK;
aTB <= "01100101100011111111110110110000";
bTB <= "11111001101001000000111011011001";
cTB <= "00100100001111010000101001111010";
dTB <= "01011110111000001100011001000000";
sel1TB <= "10010110";
sel2TB <= "00011001";
wait for T_CLK;
aTB <= "01010011110101011111101001001000";
bTB <= "10111110000001001110100011001011";
cTB <= "00000100100101110010101001001101";
dTB <= "01011000000101100110101000100101";
sel1TB <= "10101100";
sel2TB <= "10100001";
wait for T_CLK;
aTB <= "10100010101110110101101000000001";
bTB <= "11010011110011110100010111111100";
cTB <= "11111010100010010000000000111110";
dTB <= "00011011100010001101011110011010";
sel1TB <= "00111010";
sel2TB <= "10100100";
wait for T_CLK;
aTB <= "00110110011101001010100111100001";
bTB <= "01001000100010011011010001000111";
cTB <= "11000011101111000101110010101001";
dTB <= "00000001101011110011011000011111";
sel1TB <= "00110100";
sel2TB <= "01001110";
wait for T_CLK;
aTB <= "10011101110000110111110100111000";
bTB <= "00100111011000110011010000000001";
cTB <= "01011000011100000010101100100000";
dTB <= "01010011011001010100111000000011";
sel1TB <= "00100001";
sel2TB <= "11101110";
wait for T_CLK;
aTB <= "11101100111000110000011001011100";
bTB <= "01110010001110001100010000111001";
cTB <= "10010100000101101111110010001111";
dTB <= "10100011000110001100101111011111";
sel1TB <= "01111111";
sel2TB <= "00000111";
wait for T_CLK;
aTB <= "10000000100111100001111001001111";
bTB <= "10110101010111110111001110100101";
cTB <= "01010111110011010011001110011111";
dTB <= "00111111110010110101100000001111";
sel1TB <= "01011010";
sel2TB <= "11100001";
wait for T_CLK;
aTB <= "00111000010110011110001111011000";
bTB <= "01001100000011100000100110010101";
cTB <= "00111001001111000111100000101001";
dTB <= "01111101100011000100101010101000";
sel1TB <= "10101000";
sel2TB <= "10111110";
wait for T_CLK;
aTB <= "10101101010000101001010110001110";
bTB <= "00100100000001101001110100011011";
cTB <= "10101101010011110001010001101000";
dTB <= "11111000000010001100101111110010";
sel1TB <= "01111110";
sel2TB <= "00110101";
wait for T_CLK;
aTB <= "00011001101111101001101110110010";
bTB <= "00110001100101110100111111011001";
cTB <= "10010101110000001011011101010001";
dTB <= "10110111100110110101010110001001";
sel1TB <= "11100101";
sel2TB <= "00001110";
wait for T_CLK;
aTB <= "01111000010010000011000000110000";
bTB <= "00100001111000010010011110010101";
cTB <= "10011111111101111100111111001100";
dTB <= "11110010011001111000011010111111";
sel1TB <= "10000011";
sel2TB <= "11000100";
wait for T_CLK;
aTB <= "11111011010111110111111110111000";
bTB <= "10001001110110100111111011101010";
cTB <= "11110011110111010101010001011011";
dTB <= "00011000110001101001000101110010";
sel1TB <= "11100111";
sel2TB <= "10111100";
wait for T_CLK;
aTB <= "01111101111111101100000111000011";
bTB <= "00101000110111010101110110110011";
cTB <= "10011011010110101111001000111011";
dTB <= "11101100111111000010101000101111";
sel1TB <= "10010100";
sel2TB <= "10110110";
wait for T_CLK;
aTB <= "10010001110111001111000111010010";
bTB <= "01010101011000001101000110111011";
cTB <= "00001110111010101001010110001100";
dTB <= "10110110110101110000100111100010";
sel1TB <= "01110011";
sel2TB <= "01001000";
wait for T_CLK;
aTB <= "11001100001000001011011000101001";
bTB <= "11011001100000000011110110001100";
cTB <= "11010001001000101110001010011001";
dTB <= "01111110001010100010010100011111";
sel1TB <= "00101111";
sel2TB <= "00000011";
wait for T_CLK;
aTB <= "10001111011110010010010110011001";
bTB <= "01011000011000110000100010100001";
cTB <= "01011100101001010100111101011100";
dTB <= "10011000011001000011111000001000";
sel1TB <= "11101000";
sel2TB <= "11111000";
wait for T_CLK;
aTB <= "10001111000000000011011010111110";
bTB <= "00011100110001100110000011100000";
cTB <= "10001011001001111100111010001011";
dTB <= "00110001100111000100001001001011";
sel1TB <= "10100010";
sel2TB <= "01101000";
wait for T_CLK;

				
		end process uut_process;


end Behavioral;
