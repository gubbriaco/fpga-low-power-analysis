library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


package MyDefinitions is
	constant nBitsInputs : integer := 32;
	constant nBitsSels : integer := 8;
end package;